LIBRARY ieee ;
USE ieee.std_logic_1164.all ;


ENTITY transf_8bits_5bits IS
	PORT ( 	entrada : IN STD_LOGIC_VECTOR (7 downto 0) ;
				saida : OUT STD_LOGIC_VECTOR (4 DOWNTO 0)
	) ;
	END transf_8bits_5bits ;
ARCHITECTURE Behavior OF transf_8bits_5bits IS
BEGIN

	with entrada select
		saida <= "00000" when "00000000",
					"00001" when "00000001",
					"00010" when "00000010",
					"00011" when "00000011",
					"00100" when "00000100",
					"00101" when "00000101",
					"00110" when "00000110",
					"00111" when "00000111",
					"01000" when "00001000",
					"01001" when "00001001",
					"01010" when "00010000",
					"01011" when "00010001",
					"01100" when "00010010",
					"01101" when "00010011",
					"01110" when "00010100",
					"01111" when "00010101",
					"10000" when "00010110",
					"10001" when "00010111",
					"10010" when "00011000",
					"10011" when "00011001",
					"10100" when "00100000",
					"10101" when "00100001",
					"10110" when "00100010",
					"10111" when "00100011",
					"-----" when others;
END Behavior ;